
module verademo
(
	input         clk,
	input         reset,
	
	input         pal,
	input         scandouble,

	output reg    ce_pix,

	output reg    HBlank,
	output reg    HSync,
	output reg    VBlank,
	output reg    VSync,

	output  [23:0] video
);

reg   [9:0] hc;
reg   [9:0] vc;
reg   [9:0] vvc;
reg  [63:0] rnd_reg;

wire  [5:0] rnd_c = {rnd_reg[0],rnd_reg[1],rnd_reg[2],rnd_reg[2],rnd_reg[2],rnd_reg[2]};
wire [63:0] rnd;

lfsr random(rnd);

always @(posedge clk) begin
	if(scandouble) ce_pix <= 1;
		else ce_pix <= ~ce_pix;

	if(reset) begin
		hc <= 0;
		vc <= 0;
	end
	else if(ce_pix) begin
		if(hc == 637) begin
			hc <= 0;
			if(vc == (pal ? (scandouble ? 623 : 311) : (scandouble ? 523 : 261))) begin 
				vc <= 0;
				vvc <= vvc + 9'd6;
			end else begin
				vc <= vc + 1'd1;
			end
		end else begin
			hc <= hc + 1'd1;
		end

		rnd_reg <= rnd;
	end
end

always @(posedge clk) begin
	if (hc == 529) HBlank <= 1;
		else if (hc == 0) HBlank <= 0;

	if (hc == 544) begin
		HSync <= 1;

		if(pal) begin
			if(vc == (scandouble ? 609 : 304)) VSync <= 1;
				else if (vc == (scandouble ? 617 : 308)) VSync <= 0;

			if(vc == (scandouble ? 601 : 300)) VBlank <= 1;
				else if (vc == 0) VBlank <= 0;
		end
		else begin
			if(vc == (scandouble ? 490 : 245)) VSync <= 1;
				else if (vc == (scandouble ? 496 : 248)) VSync <= 0;

			if(vc == (scandouble ? 480 : 240)) VBlank <= 1;
				else if (vc == 0) VBlank <= 0;
		end
	end
	
	if (hc == 590) HSync <= 0;
end

//reg  [7:0] cos_out;
//wire [5:0] cos_g = cos_out[7:3]+6'd32;
//cos cos(vvc + {vc>>scandouble, 2'b00}, cos_out);

//assign video = (cos_g >= rnd_c) ? {cos_g - rnd_c, 2'b00} : 8'd0;

always @(posedge clk) begin
	if(pal) begin
		if(vc < (scandouble ? 400 : 200)) begin // vertical bars
			case (hc)
				0:	  video <= 24'hB4B4B4; // 75% white
				76:  video <= 24'hB4B410; // 75% yellow
				151: video <= 24'h10B4B4; // 75% cyan
				227: video <= 24'h10B410; // 75% green
				303: video <= 24'hB410B4; // 75% magenta
				379: video <= 24'hB41010; // 75% red
				454: video <= 24'h1010B4; // 75% blue
			endcase
		end
		else if (vc < (scandouble ? 467 : 233)) begin // castellations
			case (hc)
				0:	  video <= 24'h1010B4; // 75% blue
				76:  video <= 24'h101010; // 75% black
				151: video <= 24'hB410B4; // 75% magenta
				227: video <= 24'h101010; // 75% black
				303: video <= 24'h10B4B4; // 75% cyan
				379: video <= 24'h101010; // 75% black
				454: video <= 24'hB4B4B4; // 75% white
			endcase
		end
		else begin // squares
			case (hc)
				0:	  video <= 24'h10466A; // -I
				88:  video <= 24'hEBEBEB; // 100% white
				177: video <= 24'h481076; // +Q
				265: video <= 24'h101010; // 75% black
			endcase
		end
	end
	else begin // NTSC
		if(vc < (scandouble ? 320 : 160)) begin // vertical bars
			case (hc)
				0:	  video <= 24'hB4B4B4; // 75% white
				76:  video <= 24'hB4B410; // 75% yellow
				151: video <= 24'h10B4B4; // 75% cyan
				227: video <= 24'h10B410; // 75% green
				303: video <= 24'hB410B4; // 75% magenta
				379: video <= 24'hB41010; // 75% red
				454: video <= 24'h1010B4; // 75% blue
			endcase
		end
		else if (vc < (scandouble ? 373 : 187)) begin // castellations
			case (hc)
				0:	  video <= 24'h1010B4; // 75% blue
				76:  video <= 24'h101010; // 75% black
				151: video <= 24'hB410B4; // 75% magenta
				227: video <= 24'h101010; // 75% black
				303: video <= 24'h10B4B4; // 75% cyan
				379: video <= 24'h101010; // 75% black
				454: video <= 24'hB4B4B4; // 75% white
			endcase
		end
		else begin // squares
			case (hc)
				0:	  video <= 24'h10466A; // -I
				88:  video <= 24'hEBEBEB; // 100% white
				177: video <= 24'h481076; // +Q
				265: video <= 24'h101010; // 75% black
			endcase
		end
	end 

end

endmodule
